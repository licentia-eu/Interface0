/*
    Copyright (c) 2022, BogDan Vatra <bogdan@kde.org>

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <http://www.gnu.org/licenses/>.
*/
`include "Interface0_defs.v"

module Interface0(
    input ZX_CLK, /* The CK signal, sometimes referred to as PHICPU or ΦCPU is available on Lower Pin 8.
                     This clock signal is generated by the ULA and is interrupted during contended memory access.
                     On the UK 128 the ULA clock pin is connected directly to the edge connector and is inverted by TR3 to drive the Z80.
                     On the +2 the ULA clock pin is inverted by a NOT gate to generate the clock for the Z80.
                     It is then inverted again by a second NOT gate to generate the edge connector CK.
                     The CK signal is NOT connected on the Investrónica ZX Spectrum 128.
                   */

    input ZX_M1_n,  /* Machine Cycle One (output, active Low). M1, together with MREQ, indicates that the
                     current machine cycle is the op code fetch cycle of an instruction execution. M1, when
                     operating together with IORQ, indicates an interrupt acknowledge cycle.
                   */
    input ZX_MREQ_n,  /* Memory Request (output, active Low, tristate). MREQ indicates that the address
                       bus holds a valid address for a memory read or a memory write operation.
                     */

    input ZX_IORQ_n,  /* Input/Output Request (output, active Low, tristate). IORQ indicates that the lower
                       half of the address bus holds a valid I/O address for an I/O read or write operation. IORQ
                       is also generated concurrently with M1 during an interrupt acknowledge cycle to indicate
                       that an interrupt response vector can be placed on the data bus.
                     */

    input ZX_RD_n,  /* Read (output, active Low, tristate). RD indicates that the CPU wants to read data from
                     memory or an I/O device. The addressed I/O device or memory should use this signal to
                     gate data onto the CPU data bus.
                   */

    input ZX_WR_n,  /* Write (output, active Low, tristate). WR indicates that the CPU data bus contains
                     valid data to be stored at the addressed memory or I/O location
                   */

    input [15:0] ZX_ADDR, /* Address Bus (output, active High, tristate). A15-A0 form a 16-bit Address Bus,
                             which provides the addresses for memory data bus exchanges (up to 64KB) and for I/O
                             device exchanges.
                           */
    inout [7:0] ZX_DATA, /* Data Bus (input/output, active High, tristate). D7-D0 constitute an 8-bit
                            bidirectional data bus, used for data exchanges with memory and I/O
                          */

    output ZX_INT_n, /* Interrupt Request (input, active Low). An Interrupt Request is generated by I/O
                      devices. The CPU honors a request at the end of the current instruction if the internal soft-
                      ware-controlled interrupt enable flip-flop (IFF) is enabled. INT is normally wired-OR and
                      requires an external pull-up for these applications.
                    */

    output ZX_NMI, /* Nonmaskable Interrupt (input, negative edge-triggered). NMI contains a higher
                      priority than INT. NMI is always recognized at the end of the current instruction,
                      independent of the status of the interrupt enable flip-flop, and automatically forces the
                      CPU to restart at location 0066h.
                    */

    output ZX_WAIT_n, /* WAIT (input, active Low). WAIT communicates to the CPU that the addressed
                       memory or I/O devices are not ready for a data transfer. The CPU continues to enter a
                       WAIT state as long as this signal is active. Extended WAIT periods can prevent the CPU
                       from properly refreshing dynamic memory.
                     */

    output ZX_RESET_n, /* Reset (input, active Low). RESET initializes the CPU as follows: it resets the
                        interrupt enable flip-flop, clears the Program Counter and registers I and R, and sets the
                        interrupt status to Mode 0. During reset time, the address and data bus enter a
                        high-impedance state, and all control output signals enter an inactive state. RESET must be
                        active for a minimum of three full clock cycles before a reset operation is complete.
                      */

    output ZX_BUSRQ_n, /* Bus Request (input, active Low). Bus Request contains a higher priority than
                        NMI and is always recognized at the end of the current machine cycle. BUSREQ forces
                        the CPU address bus, data bus, and control signals MREQ, IORQ, RD, and WR to enter a
                        high-impedance state so that other devices can control these lines. BUSREQ is normally
                        wired OR and requires an external pull-up for these applications. Extended BUSREQ peri-
                        ods due to extensive DMA operations can prevent the CPU from properly refreshing
                        dynamic RAM.
                      */

    input ZX_BUSACK_n, /* Bus Acknowledge (output, active Low). Bus Acknowledge indicates to the
                        requesting device that the CPU address bus, data bus, and control signals MREQ, IORQ,
                        RD, and WR have entered their high-impedance states. The external circuitry can now
                        control these lines.
                      */

    // 16K/48K/128K specific
    output ZX_ROMCS, /* The ZX Spectrum 16K/48K, ZX Spectrum 128, and ZX Spectrum +2 provide ROMCS on lower pin 25.
                        By holding this pin high an external peripheral can prevent the Spectrum's ROM from driving the data bus,
                        and place its own ROM or RAM within the first 16K of the 64K memory space.
                      */

    // +2A/2B, +3/3B specific
    output ZX_ROMCS1, // All the previous models of ZX Spectrum have a single ROM chip which could be disabled to facilitate paging
    output ZX_ROMCS2, /* in external memory by pulling the ROMCS line high. The +2A/+3 and +3B however have two ROM chips and brings
                         them out to independent pins on the expansion port. The old ROMCS pin (Lower pin 25) is not used, and instead
                         Upper pin 4 and Lower pin 15 are used. These pins were both unused on the 128K, however Lower pin 15 was used
                         for composite video out on the 16K/48K.
                       */


    input ZX_DRD, // Unlike the +3, the +2A and +2B have no floppy disc controller. Amstrad's original intention was to produce an
    input ZX_DWR, // external floppy controller addon which would have connected to the expansion port on these computers.
    input ZX_MTR, /* Since the gate array is the same on all three machines, all the decoding logic is already present to generate
                     the disk read/write and motor control signals. These three signals are therefore connected through to
                     the expansion port. These signals occupy the pins which were originally used for the component video
                     signals on the 16k/48k expansion port.
                   */


    // RPi0
    input PI_MASTER_CLK,
    input SPI_CLK,
    input SPI_CS_n,
    input SPI_MOSI,
    output SPI_MISO,


    inout PI_GPIO1,
    inout PI_GPIO2,
    inout PI_GPIO3,
    inout PI_GPIO4,
    input PI_RESET
    );

reg waitData      = 1'b0;
reg romcs         = 1'b0;
reg nmi           = 1'b0;
reg resetNmi      = 1'b0;
reg haveZxData    = 1'b0;

reg [7:0] zxDataReg     = 8'd0;
reg setZxData           = 1'b0;
reg [7:0]   ioData;
reg [4:0]   bitsCounter = 5'd0;

reg sendingData         = 1'b0;
reg waitReply           = 1'b0;
reg misoData;
assign SPI_MISO = !SPI_CS_n ? misoData : 1'bz;

reg [2:0] spiClk;
always @(posedge PI_MASTER_CLK) spiClk <= {spiClk[1:0], SPI_CLK};
wire spiClkPos = (spiClk[2:1] == 2'b01);

//reg [1:0] spiClk;
//always @(posedge PI_MASTER_CLK) spiClk <= {spiClk[0], SPI_CLK};
//wire spiClkPos = (spiClk == 2'b01);

reg [2:0] zxClk;
always @(posedge PI_MASTER_CLK) zxClk <= {zxClk[1:0], ZX_CLK};
wire zxClkPos = (zxClk[2:1] == 2'b01);

reg [2:0] zxRd;
always @(posedge PI_MASTER_CLK) zxRd <= {zxRd[1:0], ZX_RD_n};
wire zxRdPos = (zxRd[2:1] == 2'b01);
wire zxRdNeg = (zxRd[2:1] == 2'b10);

wire romRead = (zxRdNeg && !ZX_MREQ_n && ~|(ZX_ADDR[15:14]));

reg [2:0] zxWr;
always @(posedge PI_MASTER_CLK) zxWr <= {zxWr[1:0], ZX_WR_n};
wire zxWrNeg = (zxWr[2:1] == 2'b10);

assign ZX_RESET_n = PI_RESET ? 0 : 1'bz;
assign ZX_ROMCS = romcs ? romcs : 1'bz;
assign ZX_WAIT_n  = !waitData;
assign ZX_NMI   = (resetNmi | nmi) ? nmi : 1'bz;
assign ZX_DATA  = setZxData ? zxDataReg : 8'bZZZZZZZZ;

assign PI_GPIO1 = romcs;
assign PI_GPIO2 = nmi;
assign PI_GPIO3 = sendingData;
assign PI_GPIO4 = haveZxData;

always @(posedge PI_MASTER_CLK) begin
  if (spiClkPos && !SPI_CS_n) begin
    misoData <= sendingData ? ioData[7] : 1'b1;
    ioData <= {ioData[6:0], SPI_MOSI};
    bitsCounter <= bitsCounter + 1;
  end

  if (bitsCounter == 5'd0 && !sendingData && !waitReply && SPI_CS_n) begin
    if (waitData) begin
      waitReply <= !ZX_RD_n;
      if (!ZX_MREQ_n) begin
        ioData <= ZX_ADDR[15:8];
      end else begin
        ioData[7] <= 1'b1;
        ioData[6] <= !ZX_RD_n;
        ioData[5] <= !ZX_WR_n;
      end
    end
    sendingData <= waitData;
  end

  if (bitsCounter == 5'd8) begin
    if (ioData[1]) begin
      romcs = ioData[7];
      if (ioData[6]) begin
        nmi <= 1'b1; // we're resetting nmi on zx clk
        resetNmi <= 1'b1;
      end
    end // if (ioData[1])

    if (sendingData) begin
      if (!ZX_MREQ_n) begin
        ioData <= ZX_ADDR[7:0];
      end else begin
        ioData <= ZX_DATA;
      end
    end else if (waitReply) begin
      haveZxData <= ioData[0];
    end

    bitsCounter <= bitsCounter + 1;
  end

  if (bitsCounter == 5'd17) begin
    if (haveZxData) begin
      zxDataReg <= ioData[7:0];
      waitData  <= 1'b0;
      setZxData <= 1'b1;
      waitReply <= 1'b0;
    end
    haveZxData  <= 1'b0;
    bitsCounter <= 5'd0;
    sendingData <= 1'b0;
  end

  if (!waitData && !setZxData) begin
    if (romRead && ZX_ADDR == `NMI_ADDR)
      romcs = 1'b1;
    if ((romRead && romcs) || ((zxRdNeg || zxWrNeg) && !ZX_IORQ_n && ZX_M1_n && ZX_ADDR == `bZX_CMD))
      waitData <= 1;
  end

  if (zxRdPos) setZxData <= 1'b0;

  if (zxClkPos) begin
    if (resetNmi) begin
      if (nmi) nmi <= 1'b0;
      else resetNmi <= 1'b0;
    end
  end // if (zxClkPos) begin

end // always @(posedge PI_MASTER_CLK) begin

endmodule
