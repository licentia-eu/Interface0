/*
    Copyright (c) 2022, BogDan Vatra <bogdan@kde.org>

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with this program.  If not, see <http://www.gnu.org/licenses/>.
*/
`include "Interface0_defs.v"

module Interface0(
    input ZX_CLK, /* The CK signal, sometimes referred to as PHICPU or ΦCPU is available on Lower Pin 8.
                     This clock signal is generated by the ULA and is interrupted during contended memory access.
                     On the UK 128 the ULA clock pin is connected directly to the edge connector and is inverted by TR3 to drive the Z80.
                     On the +2 the ULA clock pin is inverted by a NOT gate to generate the clock for the Z80.
                     It is then inverted again by a second NOT gate to generate the edge connector CK.
                     The CK signal is NOT connected on the Investrónica ZX Spectrum 128.
                   */

    input ZX_M1,  /* Machine Cycle One (output, active Low). M1, together with MREQ, indicates that the
                     current machine cycle is the op code fetch cycle of an instruction execution. M1, when
                     operating together with IORQ, indicates an interrupt acknowledge cycle.
                   */
    input ZX_MREQ,  /* Memory Request (output, active Low, tristate). MREQ indicates that the address
                       bus holds a valid address for a memory read or a memory write operation.
                     */

    input ZX_IORQ,  /* Input/Output Request (output, active Low, tristate). IORQ indicates that the lower
                       half of the address bus holds a valid I/O address for an I/O read or write operation. IORQ
                       is also generated concurrently with M1 during an interrupt acknowledge cycle to indicate
                       that an interrupt response vector can be placed on the data bus.
                     */

    input ZX_RD,  /* Read (output, active Low, tristate). RD indicates that the CPU wants to read data from
                     memory or an I/O device. The addressed I/O device or memory should use this signal to
                     gate data onto the CPU data bus.
                   */

    input ZX_WR,  /* Write (output, active Low, tristate). WR indicates that the CPU data bus contains
                     valid data to be stored at the addressed memory or I/O location
                   */

    input [15:0] ZX_ADDR, /* Address Bus (output, active High, tristate). A15-A0 form a 16-bit Address Bus,
                             which provides the addresses for memory data bus exchanges (up to 64KB) and for I/O
                             device exchanges.
                           */
    inout [7:0] ZX_DATA, /* Data Bus (input/output, active High, tristate). D7-D0 constitute an 8-bit
                            bidirectional data bus, used for data exchanges with memory and I/O
                          */

    output ZX_INT, /* Interrupt Request (input, active Low). An Interrupt Request is generated by I/O
                      devices. The CPU honors a request at the end of the current instruction if the internal soft-
                      ware-controlled interrupt enable flip-flop (IFF) is enabled. INT is normally wired-OR and
                      requires an external pull-up for these applications.
                    */

    output ZX_NMI, /* Nonmaskable Interrupt (input, negative edge-triggered). NMI contains a higher
                      priority than INT. NMI is always recognized at the end of the current instruction,
                      independent of the status of the interrupt enable flip-flop, and automatically forces the
                      CPU to restart at location 0066h.
                    */

    output ZX_WAIT, /* WAIT (input, active Low). WAIT communicates to the CPU that the addressed
                       memory or I/O devices are not ready for a data transfer. The CPU continues to enter a
                       WAIT state as long as this signal is active. Extended WAIT periods can prevent the CPU
                       from properly refreshing dynamic memory.
                     */

    output ZX_RESET, /* Reset (input, active Low). RESET initializes the CPU as follows: it resets the
                        interrupt enable flip-flop, clears the Program Counter and registers I and R, and sets the
                        interrupt status to Mode 0. During reset time, the address and data bus enter a
                        high-impedance state, and all control output signals enter an inactive state. RESET must be
                        active for a minimum of three full clock cycles before a reset operation is complete.
                      */

    output ZX_BUSRQ, /* Bus Request (input, active Low). Bus Request contains a higher priority than
                        NMI and is always recognized at the end of the current machine cycle. BUSREQ forces
                        the CPU address bus, data bus, and control signals MREQ, IORQ, RD, and WR to enter a
                        high-impedance state so that other devices can control these lines. BUSREQ is normally
                        wired OR and requires an external pull-up for these applications. Extended BUSREQ peri-
                        ods due to extensive DMA operations can prevent the CPU from properly refreshing
                        dynamic RAM.
                      */

    input ZX_BUSACK, /* Bus Acknowledge (output, active Low). Bus Acknowledge indicates to the
                        requesting device that the CPU address bus, data bus, and control signals MREQ, IORQ,
                        RD, and WR have entered their high-impedance states. The external circuitry can now
                        control these lines.
                      */

    // 16K/48K/128K specific
    output ZX_ROMCS, /* The ZX Spectrum 16K/48K, ZX Spectrum 128, and ZX Spectrum +2 provide ROMCS on lower pin 25.
                        By holding this pin high an external peripheral can prevent the Spectrum's ROM from driving the data bus,
                        and place its own ROM or RAM within the first 16K of the 64K memory space.
                      */

    // +2A/2B, +3/3B specific
    output ZX_ROMCS1, // All the previous models of ZX Spectrum have a single ROM chip which could be disabled to facilitate paging
    output ZX_ROMCS2, /* in external memory by pulling the ROMCS line high. The +2A/+3 and +3B however have two ROM chips and brings
                         them out to independent pins on the expansion port. The old ROMCS pin (Lower pin 25) is not used, and instead
                         Upper pin 4 and Lower pin 15 are used. These pins were both unused on the 128K, however Lower pin 15 was used
                         for composite video out on the 16K/48K.
                       */


    input ZX_DRD, // Unlike the +3, the +2A and +2B have no floppy disc controller. Amstrad's original intention was to produce an
    input ZX_DWR, // external floppy controller addon which would have connected to the expansion port on these computers.
    input ZX_MTR, /* Since the gate array is the same on all three machines, all the decoding logic is already present to generate
                     the disk read/write and motor control signals. These three signals are therefore connected through to
                     the expansion port. These signals occupy the pins which were originally used for the component video
                     signals on the 16k/48k expansion port.
                   */


    // RPi0
    input PI_MASTER_CLK,
    input PI_IO_CLK,
    inout PI_IO,
    input PI_MOSI,
    output PI_MISO,


    inout PI_GPIO1,
    inout PI_GPIO2,
    inout PI_GPIO3,
    inout PI_GPIO4,
    inout PI_GPIO5
    );

reg [7:0] ZX_DATA_reg = 8'd0;
reg setZxData         = 1'b0;

reg [13:0] pi_data    = 14'd0;
reg [4:0] bitsCounter = 5'd0;
reg [2:0] reset       = 3'd0;

reg piClk = 1'b0, piClkOld = 1'b0;
reg zxClk = 1'b0, zxClkOld = 1'b0;
reg m1    = 1'b0, m1Old    = 1'b0;
reg mosi  = 1'b0, mosiOld  = 1'b0;
reg miso  = 1'b0;

reg waitData  = 1'b0;
reg waitReply = 1'b0;
reg romcs     = 1'b0;
reg nmi       = 1'b0;
reg misoIoBit = 1'b0;

initial begin
  $monitor("t=%3d ZX CK=%b; M1=%b; MREQ=%b; IORQ=%b; RD=%b; WR=%b; ADDR=%b; DATA=%b; WAIT=%b; RESET=%b; ROMCS=%b, setZxData=%b",
            $time, ZX_CLK, ZX_M1, ZX_MREQ, ZX_IORQ, ZX_RD, ZX_WR, ZX_ADDR, ZX_DATA, ZX_WAIT, ZX_RESET, ZX_ROMCS, setZxData);
//
//  $monitor("t=%3d PI MASTER_CLK=%b; IO_CK=%b; IO=%b; MOSI=%b; MISO=%b; GPIO1=%b; GPIO2=%b; GPIO3=%b",
//            $time, PI_MASTER_CLK, PI_IO_CLK, PI_IO, PI_MOSI, PI_MISO, PI_GPIO1, PI_GPIO2, PI_GPIO3);
  $monitor("t=%3d IO_CK=%b; IO=%b; MOSI=%b; MISO=%b; misoIoBit=%b",
            $time, PI_IO_CLK, PI_IO, PI_MOSI, PI_MISO, misoIoBit);
end

assign ZX_ROMCS = ~|romcs;
assign ZX_WAIT  = ~|waitData;
assign ZX_RESET = ~|reset;
assign ZX_NMI   = ~|nmi;
assign ZX_DATA  = (!ZX_RD && setZxData) ? ZX_DATA_reg : 8'bZZZZZZZZ;

assign PI_MISO = miso;
assign PI_IO   = !PI_MOSI ? misoIoBit : 1'bz;

always @(posedge PI_MASTER_CLK) begin
  zxClkOld <= ZX_CLK;
  zxClk <= zxClkOld;
  if (zxClk == 1'b0 && zxClkOld == 1'b1) begin // zx_clk pos edge
    if (nmi) begin
      m1Old <= ZX_M1;
      m1 <= m1Old;
      if (m1 == 0 && m1Old == 1) nmi <= 0;// wait untill we have an M1 neg edge
    end

    if (setZxData && ZX_RD) setZxData <= 0;
    if (|reset) reset <= reset - 1;

    if (!waitData && !setZxData) begin
      if (!ZX_ROMCS && !ZX_MREQ && !ZX_RD && ZX_ADDR[15:14] == 2'b00) begin
        bitsCounter <= 5'd13;
        waitData <= 1;
        pi_data <= ZX_ADDR[13:0];
        miso <= 1; // what will happen if we're in a middle of a MOSI?
        waitReply <= 1'b1;
      end

      if (!ZX_IORQ && (!ZX_RD || !ZX_WR)) begin
        if (ZX_ADDR == `bZX_CMD) begin
          pi_data[13:5] <= {!ZX_RD, ZX_DATA};
          waitData <= !ZX_RD;
          waitReply <= !ZX_WR;
          bitsCounter <= 5'd9;
          miso <= 1; // what will happen if we're in a middle of a MOSI?
        end
      end
    end // if (!waitData) begin
  end // if (zxClk == 1'b1 && zxClkOld == 1'b0) begin



  piClkOld <= PI_IO_CLK;
  piClk <= piClkOld;
  if (piClk == 1'b0 && piClkOld == 1'b1) begin // pi_clk pos edge
    if (PI_MOSI) begin // read from PI
      pi_data <= {pi_data[12:0], PI_IO};
      bitsCounter <= bitsCounter + 1;
    end else begin // send to PI
      bitsCounter <= bitsCounter - 1;
      misoIoBit <= pi_data[13];
      pi_data <= {pi_data[12:0], 1'b0};
      if (~|bitsCounter) begin
        miso <= 0;
        if (!waitReply) begin
          waitData <= 0;
        end
      end
    end
  end // if (piClk == 1'b1 && piClkOld == 1'b0) begin



  mosiOld <= PI_MOSI;
  mosi <= mosiOld;
  if (mosi == 1'b0 && mosiOld == 1'b1) begin// mosi pos edge
    bitsCounter <= 0;
  end else if (mosi == 1'b1 && mosiOld == 1'b0) begin // mosi neg edge
    waitReply <= 1'b0;
    if (bitsCounter == 5'd4) begin // simple command
      if (~|(pi_data[3:0] & `CMDS)) begin
        romcs <= |(pi_data[3:0] & `ROMCS_CMD);
        reset <= (|(pi_data[3:0] & `RESET_CMD)) ? `RESET_COUNT : 3'd0;
        nmi <= |(pi_data[3:0] & `NMI_CMD);
      end
    end else begin
      if (waitData && bitsCounter == 5'd8) begin
        ZX_DATA_reg <= pi_data[7:0];
        setZxData <= 1;
        waitData <= 0;
      end
    end
  end // else if (mosi == 1'b0 && mosiOld == 1'b1) begin
end

endmodule
